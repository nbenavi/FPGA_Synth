module Addcout18 (input [17:0] I0, input [17:0] I1, output [17:0] O, output  COUT);
wire  inst0_O;
wire  inst1_CO;
wire  inst2_O;
wire  inst3_CO;
wire  inst4_O;
wire  inst5_CO;
wire  inst6_O;
wire  inst7_CO;
wire  inst8_O;
wire  inst9_CO;
wire  inst10_O;
wire  inst11_CO;
wire  inst12_O;
wire  inst13_CO;
wire  inst14_O;
wire  inst15_CO;
wire  inst16_O;
wire  inst17_CO;
wire  inst18_O;
wire  inst19_CO;
wire  inst20_O;
wire  inst21_CO;
wire  inst22_O;
wire  inst23_CO;
wire  inst24_O;
wire  inst25_CO;
wire  inst26_O;
wire  inst27_CO;
wire  inst28_O;
wire  inst29_CO;
wire  inst30_O;
wire  inst31_CO;
wire  inst32_O;
wire  inst33_CO;
wire  inst34_O;
wire  inst35_CO;
SB_LUT4 #(.LUT_INIT(16'hC33C)) inst0 (.I0(1'b0), .I1(I0[0]), .I2(I1[0]), .I3(1'b0), .O(inst0_O));
SB_CARRY inst1 (.I0(I0[0]), .I1(I1[0]), .CI(1'b0), .CO(inst1_CO));
SB_LUT4 #(.LUT_INIT(16'hC33C)) inst2 (.I0(1'b0), .I1(I0[1]), .I2(I1[1]), .I3(inst1_CO), .O(inst2_O));
SB_CARRY inst3 (.I0(I0[1]), .I1(I1[1]), .CI(inst1_CO), .CO(inst3_CO));
SB_LUT4 #(.LUT_INIT(16'hC33C)) inst4 (.I0(1'b0), .I1(I0[2]), .I2(I1[2]), .I3(inst3_CO), .O(inst4_O));
SB_CARRY inst5 (.I0(I0[2]), .I1(I1[2]), .CI(inst3_CO), .CO(inst5_CO));
SB_LUT4 #(.LUT_INIT(16'hC33C)) inst6 (.I0(1'b0), .I1(I0[3]), .I2(I1[3]), .I3(inst5_CO), .O(inst6_O));
SB_CARRY inst7 (.I0(I0[3]), .I1(I1[3]), .CI(inst5_CO), .CO(inst7_CO));
SB_LUT4 #(.LUT_INIT(16'hC33C)) inst8 (.I0(1'b0), .I1(I0[4]), .I2(I1[4]), .I3(inst7_CO), .O(inst8_O));
SB_CARRY inst9 (.I0(I0[4]), .I1(I1[4]), .CI(inst7_CO), .CO(inst9_CO));
SB_LUT4 #(.LUT_INIT(16'hC33C)) inst10 (.I0(1'b0), .I1(I0[5]), .I2(I1[5]), .I3(inst9_CO), .O(inst10_O));
SB_CARRY inst11 (.I0(I0[5]), .I1(I1[5]), .CI(inst9_CO), .CO(inst11_CO));
SB_LUT4 #(.LUT_INIT(16'hC33C)) inst12 (.I0(1'b0), .I1(I0[6]), .I2(I1[6]), .I3(inst11_CO), .O(inst12_O));
SB_CARRY inst13 (.I0(I0[6]), .I1(I1[6]), .CI(inst11_CO), .CO(inst13_CO));
SB_LUT4 #(.LUT_INIT(16'hC33C)) inst14 (.I0(1'b0), .I1(I0[7]), .I2(I1[7]), .I3(inst13_CO), .O(inst14_O));
SB_CARRY inst15 (.I0(I0[7]), .I1(I1[7]), .CI(inst13_CO), .CO(inst15_CO));
SB_LUT4 #(.LUT_INIT(16'hC33C)) inst16 (.I0(1'b0), .I1(I0[8]), .I2(I1[8]), .I3(inst15_CO), .O(inst16_O));
SB_CARRY inst17 (.I0(I0[8]), .I1(I1[8]), .CI(inst15_CO), .CO(inst17_CO));
SB_LUT4 #(.LUT_INIT(16'hC33C)) inst18 (.I0(1'b0), .I1(I0[9]), .I2(I1[9]), .I3(inst17_CO), .O(inst18_O));
SB_CARRY inst19 (.I0(I0[9]), .I1(I1[9]), .CI(inst17_CO), .CO(inst19_CO));
SB_LUT4 #(.LUT_INIT(16'hC33C)) inst20 (.I0(1'b0), .I1(I0[10]), .I2(I1[10]), .I3(inst19_CO), .O(inst20_O));
SB_CARRY inst21 (.I0(I0[10]), .I1(I1[10]), .CI(inst19_CO), .CO(inst21_CO));
SB_LUT4 #(.LUT_INIT(16'hC33C)) inst22 (.I0(1'b0), .I1(I0[11]), .I2(I1[11]), .I3(inst21_CO), .O(inst22_O));
SB_CARRY inst23 (.I0(I0[11]), .I1(I1[11]), .CI(inst21_CO), .CO(inst23_CO));
SB_LUT4 #(.LUT_INIT(16'hC33C)) inst24 (.I0(1'b0), .I1(I0[12]), .I2(I1[12]), .I3(inst23_CO), .O(inst24_O));
SB_CARRY inst25 (.I0(I0[12]), .I1(I1[12]), .CI(inst23_CO), .CO(inst25_CO));
SB_LUT4 #(.LUT_INIT(16'hC33C)) inst26 (.I0(1'b0), .I1(I0[13]), .I2(I1[13]), .I3(inst25_CO), .O(inst26_O));
SB_CARRY inst27 (.I0(I0[13]), .I1(I1[13]), .CI(inst25_CO), .CO(inst27_CO));
SB_LUT4 #(.LUT_INIT(16'hC33C)) inst28 (.I0(1'b0), .I1(I0[14]), .I2(I1[14]), .I3(inst27_CO), .O(inst28_O));
SB_CARRY inst29 (.I0(I0[14]), .I1(I1[14]), .CI(inst27_CO), .CO(inst29_CO));
SB_LUT4 #(.LUT_INIT(16'hC33C)) inst30 (.I0(1'b0), .I1(I0[15]), .I2(I1[15]), .I3(inst29_CO), .O(inst30_O));
SB_CARRY inst31 (.I0(I0[15]), .I1(I1[15]), .CI(inst29_CO), .CO(inst31_CO));
SB_LUT4 #(.LUT_INIT(16'hC33C)) inst32 (.I0(1'b0), .I1(I0[16]), .I2(I1[16]), .I3(inst31_CO), .O(inst32_O));
SB_CARRY inst33 (.I0(I0[16]), .I1(I1[16]), .CI(inst31_CO), .CO(inst33_CO));
SB_LUT4 #(.LUT_INIT(16'hC33C)) inst34 (.I0(1'b0), .I1(I0[17]), .I2(I1[17]), .I3(inst33_CO), .O(inst34_O));
SB_CARRY inst35 (.I0(I0[17]), .I1(I1[17]), .CI(inst33_CO), .CO(inst35_CO));
assign O = {inst34_O,inst32_O,inst30_O,inst28_O,inst26_O,inst24_O,inst22_O,inst20_O,inst18_O,inst16_O,inst14_O,inst12_O,inst10_O,inst8_O,inst6_O,inst4_O,inst2_O,inst0_O};
assign COUT = inst35_CO;
endmodule

module Register18 (input [17:0] I, output [17:0] O, input  CLK);
wire  inst0_Q;
wire  inst1_Q;
wire  inst2_Q;
wire  inst3_Q;
wire  inst4_Q;
wire  inst5_Q;
wire  inst6_Q;
wire  inst7_Q;
wire  inst8_Q;
wire  inst9_Q;
wire  inst10_Q;
wire  inst11_Q;
wire  inst12_Q;
wire  inst13_Q;
wire  inst14_Q;
wire  inst15_Q;
wire  inst16_Q;
wire  inst17_Q;
SB_DFF inst0 (.C(CLK), .D(I[0]), .Q(inst0_Q));
SB_DFF inst1 (.C(CLK), .D(I[1]), .Q(inst1_Q));
SB_DFF inst2 (.C(CLK), .D(I[2]), .Q(inst2_Q));
SB_DFF inst3 (.C(CLK), .D(I[3]), .Q(inst3_Q));
SB_DFF inst4 (.C(CLK), .D(I[4]), .Q(inst4_Q));
SB_DFF inst5 (.C(CLK), .D(I[5]), .Q(inst5_Q));
SB_DFF inst6 (.C(CLK), .D(I[6]), .Q(inst6_Q));
SB_DFF inst7 (.C(CLK), .D(I[7]), .Q(inst7_Q));
SB_DFF inst8 (.C(CLK), .D(I[8]), .Q(inst8_Q));
SB_DFF inst9 (.C(CLK), .D(I[9]), .Q(inst9_Q));
SB_DFF inst10 (.C(CLK), .D(I[10]), .Q(inst10_Q));
SB_DFF inst11 (.C(CLK), .D(I[11]), .Q(inst11_Q));
SB_DFF inst12 (.C(CLK), .D(I[12]), .Q(inst12_Q));
SB_DFF inst13 (.C(CLK), .D(I[13]), .Q(inst13_Q));
SB_DFF inst14 (.C(CLK), .D(I[14]), .Q(inst14_Q));
SB_DFF inst15 (.C(CLK), .D(I[15]), .Q(inst15_Q));
SB_DFF inst16 (.C(CLK), .D(I[16]), .Q(inst16_Q));
SB_DFF inst17 (.C(CLK), .D(I[17]), .Q(inst17_Q));
assign O = {inst17_Q,inst16_Q,inst15_Q,inst14_Q,inst13_Q,inst12_Q,inst11_Q,inst10_Q,inst9_Q,inst8_Q,inst7_Q,inst6_Q,inst5_Q,inst4_Q,inst3_Q,inst2_Q,inst1_Q,inst0_Q};
endmodule

module Counter18 (output [17:0] O, output  COUT, input  CLK);
wire [17:0] inst0_O;
wire  inst0_COUT;
wire [17:0] inst1_O;
Addcout18 inst0 (.I0(inst1_O), .I1({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1}), .O(inst0_O), .COUT(inst0_COUT));
Register18 inst1 (.I(inst0_O), .O(inst1_O), .CLK(CLK));
assign O = inst1_O;
assign COUT = inst0_COUT;
endmodule

module Addcout27 (input [26:0] I0, input [26:0] I1, output [26:0] O, output  COUT);
wire  inst0_O;
wire  inst1_CO;
wire  inst2_O;
wire  inst3_CO;
wire  inst4_O;
wire  inst5_CO;
wire  inst6_O;
wire  inst7_CO;
wire  inst8_O;
wire  inst9_CO;
wire  inst10_O;
wire  inst11_CO;
wire  inst12_O;
wire  inst13_CO;
wire  inst14_O;
wire  inst15_CO;
wire  inst16_O;
wire  inst17_CO;
wire  inst18_O;
wire  inst19_CO;
wire  inst20_O;
wire  inst21_CO;
wire  inst22_O;
wire  inst23_CO;
wire  inst24_O;
wire  inst25_CO;
wire  inst26_O;
wire  inst27_CO;
wire  inst28_O;
wire  inst29_CO;
wire  inst30_O;
wire  inst31_CO;
wire  inst32_O;
wire  inst33_CO;
wire  inst34_O;
wire  inst35_CO;
wire  inst36_O;
wire  inst37_CO;
wire  inst38_O;
wire  inst39_CO;
wire  inst40_O;
wire  inst41_CO;
wire  inst42_O;
wire  inst43_CO;
wire  inst44_O;
wire  inst45_CO;
wire  inst46_O;
wire  inst47_CO;
wire  inst48_O;
wire  inst49_CO;
wire  inst50_O;
wire  inst51_CO;
wire  inst52_O;
wire  inst53_CO;
SB_LUT4 #(.LUT_INIT(16'hC33C)) inst0 (.I0(1'b0), .I1(I0[0]), .I2(I1[0]), .I3(1'b0), .O(inst0_O));
SB_CARRY inst1 (.I0(I0[0]), .I1(I1[0]), .CI(1'b0), .CO(inst1_CO));
SB_LUT4 #(.LUT_INIT(16'hC33C)) inst2 (.I0(1'b0), .I1(I0[1]), .I2(I1[1]), .I3(inst1_CO), .O(inst2_O));
SB_CARRY inst3 (.I0(I0[1]), .I1(I1[1]), .CI(inst1_CO), .CO(inst3_CO));
SB_LUT4 #(.LUT_INIT(16'hC33C)) inst4 (.I0(1'b0), .I1(I0[2]), .I2(I1[2]), .I3(inst3_CO), .O(inst4_O));
SB_CARRY inst5 (.I0(I0[2]), .I1(I1[2]), .CI(inst3_CO), .CO(inst5_CO));
SB_LUT4 #(.LUT_INIT(16'hC33C)) inst6 (.I0(1'b0), .I1(I0[3]), .I2(I1[3]), .I3(inst5_CO), .O(inst6_O));
SB_CARRY inst7 (.I0(I0[3]), .I1(I1[3]), .CI(inst5_CO), .CO(inst7_CO));
SB_LUT4 #(.LUT_INIT(16'hC33C)) inst8 (.I0(1'b0), .I1(I0[4]), .I2(I1[4]), .I3(inst7_CO), .O(inst8_O));
SB_CARRY inst9 (.I0(I0[4]), .I1(I1[4]), .CI(inst7_CO), .CO(inst9_CO));
SB_LUT4 #(.LUT_INIT(16'hC33C)) inst10 (.I0(1'b0), .I1(I0[5]), .I2(I1[5]), .I3(inst9_CO), .O(inst10_O));
SB_CARRY inst11 (.I0(I0[5]), .I1(I1[5]), .CI(inst9_CO), .CO(inst11_CO));
SB_LUT4 #(.LUT_INIT(16'hC33C)) inst12 (.I0(1'b0), .I1(I0[6]), .I2(I1[6]), .I3(inst11_CO), .O(inst12_O));
SB_CARRY inst13 (.I0(I0[6]), .I1(I1[6]), .CI(inst11_CO), .CO(inst13_CO));
SB_LUT4 #(.LUT_INIT(16'hC33C)) inst14 (.I0(1'b0), .I1(I0[7]), .I2(I1[7]), .I3(inst13_CO), .O(inst14_O));
SB_CARRY inst15 (.I0(I0[7]), .I1(I1[7]), .CI(inst13_CO), .CO(inst15_CO));
SB_LUT4 #(.LUT_INIT(16'hC33C)) inst16 (.I0(1'b0), .I1(I0[8]), .I2(I1[8]), .I3(inst15_CO), .O(inst16_O));
SB_CARRY inst17 (.I0(I0[8]), .I1(I1[8]), .CI(inst15_CO), .CO(inst17_CO));
SB_LUT4 #(.LUT_INIT(16'hC33C)) inst18 (.I0(1'b0), .I1(I0[9]), .I2(I1[9]), .I3(inst17_CO), .O(inst18_O));
SB_CARRY inst19 (.I0(I0[9]), .I1(I1[9]), .CI(inst17_CO), .CO(inst19_CO));
SB_LUT4 #(.LUT_INIT(16'hC33C)) inst20 (.I0(1'b0), .I1(I0[10]), .I2(I1[10]), .I3(inst19_CO), .O(inst20_O));
SB_CARRY inst21 (.I0(I0[10]), .I1(I1[10]), .CI(inst19_CO), .CO(inst21_CO));
SB_LUT4 #(.LUT_INIT(16'hC33C)) inst22 (.I0(1'b0), .I1(I0[11]), .I2(I1[11]), .I3(inst21_CO), .O(inst22_O));
SB_CARRY inst23 (.I0(I0[11]), .I1(I1[11]), .CI(inst21_CO), .CO(inst23_CO));
SB_LUT4 #(.LUT_INIT(16'hC33C)) inst24 (.I0(1'b0), .I1(I0[12]), .I2(I1[12]), .I3(inst23_CO), .O(inst24_O));
SB_CARRY inst25 (.I0(I0[12]), .I1(I1[12]), .CI(inst23_CO), .CO(inst25_CO));
SB_LUT4 #(.LUT_INIT(16'hC33C)) inst26 (.I0(1'b0), .I1(I0[13]), .I2(I1[13]), .I3(inst25_CO), .O(inst26_O));
SB_CARRY inst27 (.I0(I0[13]), .I1(I1[13]), .CI(inst25_CO), .CO(inst27_CO));
SB_LUT4 #(.LUT_INIT(16'hC33C)) inst28 (.I0(1'b0), .I1(I0[14]), .I2(I1[14]), .I3(inst27_CO), .O(inst28_O));
SB_CARRY inst29 (.I0(I0[14]), .I1(I1[14]), .CI(inst27_CO), .CO(inst29_CO));
SB_LUT4 #(.LUT_INIT(16'hC33C)) inst30 (.I0(1'b0), .I1(I0[15]), .I2(I1[15]), .I3(inst29_CO), .O(inst30_O));
SB_CARRY inst31 (.I0(I0[15]), .I1(I1[15]), .CI(inst29_CO), .CO(inst31_CO));
SB_LUT4 #(.LUT_INIT(16'hC33C)) inst32 (.I0(1'b0), .I1(I0[16]), .I2(I1[16]), .I3(inst31_CO), .O(inst32_O));
SB_CARRY inst33 (.I0(I0[16]), .I1(I1[16]), .CI(inst31_CO), .CO(inst33_CO));
SB_LUT4 #(.LUT_INIT(16'hC33C)) inst34 (.I0(1'b0), .I1(I0[17]), .I2(I1[17]), .I3(inst33_CO), .O(inst34_O));
SB_CARRY inst35 (.I0(I0[17]), .I1(I1[17]), .CI(inst33_CO), .CO(inst35_CO));
SB_LUT4 #(.LUT_INIT(16'hC33C)) inst36 (.I0(1'b0), .I1(I0[18]), .I2(I1[18]), .I3(inst35_CO), .O(inst36_O));
SB_CARRY inst37 (.I0(I0[18]), .I1(I1[18]), .CI(inst35_CO), .CO(inst37_CO));
SB_LUT4 #(.LUT_INIT(16'hC33C)) inst38 (.I0(1'b0), .I1(I0[19]), .I2(I1[19]), .I3(inst37_CO), .O(inst38_O));
SB_CARRY inst39 (.I0(I0[19]), .I1(I1[19]), .CI(inst37_CO), .CO(inst39_CO));
SB_LUT4 #(.LUT_INIT(16'hC33C)) inst40 (.I0(1'b0), .I1(I0[20]), .I2(I1[20]), .I3(inst39_CO), .O(inst40_O));
SB_CARRY inst41 (.I0(I0[20]), .I1(I1[20]), .CI(inst39_CO), .CO(inst41_CO));
SB_LUT4 #(.LUT_INIT(16'hC33C)) inst42 (.I0(1'b0), .I1(I0[21]), .I2(I1[21]), .I3(inst41_CO), .O(inst42_O));
SB_CARRY inst43 (.I0(I0[21]), .I1(I1[21]), .CI(inst41_CO), .CO(inst43_CO));
SB_LUT4 #(.LUT_INIT(16'hC33C)) inst44 (.I0(1'b0), .I1(I0[22]), .I2(I1[22]), .I3(inst43_CO), .O(inst44_O));
SB_CARRY inst45 (.I0(I0[22]), .I1(I1[22]), .CI(inst43_CO), .CO(inst45_CO));
SB_LUT4 #(.LUT_INIT(16'hC33C)) inst46 (.I0(1'b0), .I1(I0[23]), .I2(I1[23]), .I3(inst45_CO), .O(inst46_O));
SB_CARRY inst47 (.I0(I0[23]), .I1(I1[23]), .CI(inst45_CO), .CO(inst47_CO));
SB_LUT4 #(.LUT_INIT(16'hC33C)) inst48 (.I0(1'b0), .I1(I0[24]), .I2(I1[24]), .I3(inst47_CO), .O(inst48_O));
SB_CARRY inst49 (.I0(I0[24]), .I1(I1[24]), .CI(inst47_CO), .CO(inst49_CO));
SB_LUT4 #(.LUT_INIT(16'hC33C)) inst50 (.I0(1'b0), .I1(I0[25]), .I2(I1[25]), .I3(inst49_CO), .O(inst50_O));
SB_CARRY inst51 (.I0(I0[25]), .I1(I1[25]), .CI(inst49_CO), .CO(inst51_CO));
SB_LUT4 #(.LUT_INIT(16'hC33C)) inst52 (.I0(1'b0), .I1(I0[26]), .I2(I1[26]), .I3(inst51_CO), .O(inst52_O));
SB_CARRY inst53 (.I0(I0[26]), .I1(I1[26]), .CI(inst51_CO), .CO(inst53_CO));
assign O = {inst52_O,inst50_O,inst48_O,inst46_O,inst44_O,inst42_O,inst40_O,inst38_O,inst36_O,inst34_O,inst32_O,inst30_O,inst28_O,inst26_O,inst24_O,inst22_O,inst20_O,inst18_O,inst16_O,inst14_O,inst12_O,inst10_O,inst8_O,inst6_O,inst4_O,inst2_O,inst0_O};
assign COUT = inst53_CO;
endmodule

module Register27 (input [26:0] I, output [26:0] O, input  CLK);
wire  inst0_Q;
wire  inst1_Q;
wire  inst2_Q;
wire  inst3_Q;
wire  inst4_Q;
wire  inst5_Q;
wire  inst6_Q;
wire  inst7_Q;
wire  inst8_Q;
wire  inst9_Q;
wire  inst10_Q;
wire  inst11_Q;
wire  inst12_Q;
wire  inst13_Q;
wire  inst14_Q;
wire  inst15_Q;
wire  inst16_Q;
wire  inst17_Q;
wire  inst18_Q;
wire  inst19_Q;
wire  inst20_Q;
wire  inst21_Q;
wire  inst22_Q;
wire  inst23_Q;
wire  inst24_Q;
wire  inst25_Q;
wire  inst26_Q;
SB_DFF inst0 (.C(CLK), .D(I[0]), .Q(inst0_Q));
SB_DFF inst1 (.C(CLK), .D(I[1]), .Q(inst1_Q));
SB_DFF inst2 (.C(CLK), .D(I[2]), .Q(inst2_Q));
SB_DFF inst3 (.C(CLK), .D(I[3]), .Q(inst3_Q));
SB_DFF inst4 (.C(CLK), .D(I[4]), .Q(inst4_Q));
SB_DFF inst5 (.C(CLK), .D(I[5]), .Q(inst5_Q));
SB_DFF inst6 (.C(CLK), .D(I[6]), .Q(inst6_Q));
SB_DFF inst7 (.C(CLK), .D(I[7]), .Q(inst7_Q));
SB_DFF inst8 (.C(CLK), .D(I[8]), .Q(inst8_Q));
SB_DFF inst9 (.C(CLK), .D(I[9]), .Q(inst9_Q));
SB_DFF inst10 (.C(CLK), .D(I[10]), .Q(inst10_Q));
SB_DFF inst11 (.C(CLK), .D(I[11]), .Q(inst11_Q));
SB_DFF inst12 (.C(CLK), .D(I[12]), .Q(inst12_Q));
SB_DFF inst13 (.C(CLK), .D(I[13]), .Q(inst13_Q));
SB_DFF inst14 (.C(CLK), .D(I[14]), .Q(inst14_Q));
SB_DFF inst15 (.C(CLK), .D(I[15]), .Q(inst15_Q));
SB_DFF inst16 (.C(CLK), .D(I[16]), .Q(inst16_Q));
SB_DFF inst17 (.C(CLK), .D(I[17]), .Q(inst17_Q));
SB_DFF inst18 (.C(CLK), .D(I[18]), .Q(inst18_Q));
SB_DFF inst19 (.C(CLK), .D(I[19]), .Q(inst19_Q));
SB_DFF inst20 (.C(CLK), .D(I[20]), .Q(inst20_Q));
SB_DFF inst21 (.C(CLK), .D(I[21]), .Q(inst21_Q));
SB_DFF inst22 (.C(CLK), .D(I[22]), .Q(inst22_Q));
SB_DFF inst23 (.C(CLK), .D(I[23]), .Q(inst23_Q));
SB_DFF inst24 (.C(CLK), .D(I[24]), .Q(inst24_Q));
SB_DFF inst25 (.C(CLK), .D(I[25]), .Q(inst25_Q));
SB_DFF inst26 (.C(CLK), .D(I[26]), .Q(inst26_Q));
assign O = {inst26_Q,inst25_Q,inst24_Q,inst23_Q,inst22_Q,inst21_Q,inst20_Q,inst19_Q,inst18_Q,inst17_Q,inst16_Q,inst15_Q,inst14_Q,inst13_Q,inst12_Q,inst11_Q,inst10_Q,inst9_Q,inst8_Q,inst7_Q,inst6_Q,inst5_Q,inst4_Q,inst3_Q,inst2_Q,inst1_Q,inst0_Q};
endmodule

module Counter27 (output [26:0] O, output  COUT, input  CLK);
wire [26:0] inst0_O;
wire  inst0_COUT;
wire [26:0] inst1_O;
Addcout27 inst0 (.I0(inst1_O), .I1({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1}), .O(inst0_O), .COUT(inst0_COUT));
Register27 inst1 (.I(inst0_O), .O(inst1_O), .CLK(CLK));
assign O = inst1_O;
assign COUT = inst0_COUT;
endmodule

module Addcout2 (input [1:0] I0, input [1:0] I1, output [1:0] O, output  COUT);
wire  inst0_O;
wire  inst1_CO;
wire  inst2_O;
wire  inst3_CO;
SB_LUT4 #(.LUT_INIT(16'hC33C)) inst0 (.I0(1'b0), .I1(I0[0]), .I2(I1[0]), .I3(1'b0), .O(inst0_O));
SB_CARRY inst1 (.I0(I0[0]), .I1(I1[0]), .CI(1'b0), .CO(inst1_CO));
SB_LUT4 #(.LUT_INIT(16'hC33C)) inst2 (.I0(1'b0), .I1(I0[1]), .I2(I1[1]), .I3(inst1_CO), .O(inst2_O));
SB_CARRY inst3 (.I0(I0[1]), .I1(I1[1]), .CI(inst1_CO), .CO(inst3_CO));
assign O = {inst2_O,inst0_O};
assign COUT = inst3_CO;
endmodule

module Register2CE (input [1:0] I, output [1:0] O, input  CLK, input  CE);
wire  inst0_Q;
wire  inst1_Q;
SB_DFFE inst0 (.C(CLK), .E(CE), .D(I[0]), .Q(inst0_Q));
SB_DFFE inst1 (.C(CLK), .E(CE), .D(I[1]), .Q(inst1_Q));
assign O = {inst1_Q,inst0_Q};
endmodule

module Counter2CE (output [1:0] O, output  COUT, input  CLK, input  CE);
wire [1:0] inst0_O;
wire  inst0_COUT;
wire [1:0] inst1_O;
Addcout2 inst0 (.I0(inst1_O), .I1({1'b0,1'b1}), .O(inst0_O), .COUT(inst0_COUT));
Register2CE inst1 (.I(inst0_O), .O(inst1_O), .CLK(CLK), .CE(CE));
assign O = inst1_O;
assign COUT = inst0_COUT;
endmodule

module Addcout8 (input [7:0] I0, input [7:0] I1, output [7:0] O, output  COUT);
wire  inst0_O;
wire  inst1_CO;
wire  inst2_O;
wire  inst3_CO;
wire  inst4_O;
wire  inst5_CO;
wire  inst6_O;
wire  inst7_CO;
wire  inst8_O;
wire  inst9_CO;
wire  inst10_O;
wire  inst11_CO;
wire  inst12_O;
wire  inst13_CO;
wire  inst14_O;
wire  inst15_CO;
SB_LUT4 #(.LUT_INIT(16'hC33C)) inst0 (.I0(1'b0), .I1(I0[0]), .I2(I1[0]), .I3(1'b0), .O(inst0_O));
SB_CARRY inst1 (.I0(I0[0]), .I1(I1[0]), .CI(1'b0), .CO(inst1_CO));
SB_LUT4 #(.LUT_INIT(16'hC33C)) inst2 (.I0(1'b0), .I1(I0[1]), .I2(I1[1]), .I3(inst1_CO), .O(inst2_O));
SB_CARRY inst3 (.I0(I0[1]), .I1(I1[1]), .CI(inst1_CO), .CO(inst3_CO));
SB_LUT4 #(.LUT_INIT(16'hC33C)) inst4 (.I0(1'b0), .I1(I0[2]), .I2(I1[2]), .I3(inst3_CO), .O(inst4_O));
SB_CARRY inst5 (.I0(I0[2]), .I1(I1[2]), .CI(inst3_CO), .CO(inst5_CO));
SB_LUT4 #(.LUT_INIT(16'hC33C)) inst6 (.I0(1'b0), .I1(I0[3]), .I2(I1[3]), .I3(inst5_CO), .O(inst6_O));
SB_CARRY inst7 (.I0(I0[3]), .I1(I1[3]), .CI(inst5_CO), .CO(inst7_CO));
SB_LUT4 #(.LUT_INIT(16'hC33C)) inst8 (.I0(1'b0), .I1(I0[4]), .I2(I1[4]), .I3(inst7_CO), .O(inst8_O));
SB_CARRY inst9 (.I0(I0[4]), .I1(I1[4]), .CI(inst7_CO), .CO(inst9_CO));
SB_LUT4 #(.LUT_INIT(16'hC33C)) inst10 (.I0(1'b0), .I1(I0[5]), .I2(I1[5]), .I3(inst9_CO), .O(inst10_O));
SB_CARRY inst11 (.I0(I0[5]), .I1(I1[5]), .CI(inst9_CO), .CO(inst11_CO));
SB_LUT4 #(.LUT_INIT(16'hC33C)) inst12 (.I0(1'b0), .I1(I0[6]), .I2(I1[6]), .I3(inst11_CO), .O(inst12_O));
SB_CARRY inst13 (.I0(I0[6]), .I1(I1[6]), .CI(inst11_CO), .CO(inst13_CO));
SB_LUT4 #(.LUT_INIT(16'hC33C)) inst14 (.I0(1'b0), .I1(I0[7]), .I2(I1[7]), .I3(inst13_CO), .O(inst14_O));
SB_CARRY inst15 (.I0(I0[7]), .I1(I1[7]), .CI(inst13_CO), .CO(inst15_CO));
assign O = {inst14_O,inst12_O,inst10_O,inst8_O,inst6_O,inst4_O,inst2_O,inst0_O};
assign COUT = inst15_CO;
endmodule

module Register8 (input [7:0] I, output [7:0] O, input  CLK);
wire  inst0_Q;
wire  inst1_Q;
wire  inst2_Q;
wire  inst3_Q;
wire  inst4_Q;
wire  inst5_Q;
wire  inst6_Q;
wire  inst7_Q;
SB_DFF inst0 (.C(CLK), .D(I[0]), .Q(inst0_Q));
SB_DFF inst1 (.C(CLK), .D(I[1]), .Q(inst1_Q));
SB_DFF inst2 (.C(CLK), .D(I[2]), .Q(inst2_Q));
SB_DFF inst3 (.C(CLK), .D(I[3]), .Q(inst3_Q));
SB_DFF inst4 (.C(CLK), .D(I[4]), .Q(inst4_Q));
SB_DFF inst5 (.C(CLK), .D(I[5]), .Q(inst5_Q));
SB_DFF inst6 (.C(CLK), .D(I[6]), .Q(inst6_Q));
SB_DFF inst7 (.C(CLK), .D(I[7]), .Q(inst7_Q));
assign O = {inst7_Q,inst6_Q,inst5_Q,inst4_Q,inst3_Q,inst2_Q,inst1_Q,inst0_Q};
endmodule

module Counter8 (output [7:0] O, output  COUT, input  CLK);
wire [7:0] inst0_O;
wire  inst0_COUT;
wire [7:0] inst1_O;
Addcout8 inst0 (.I0(inst1_O), .I1({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1}), .O(inst0_O), .COUT(inst0_COUT));
Register8 inst1 (.I(inst0_O), .O(inst1_O), .CLK(CLK));
assign O = inst1_O;
assign COUT = inst0_COUT;
endmodule

module Addcincout5 (input [4:0] I0, input [4:0] I1, input  CIN, output [4:0] O, output  COUT);
wire  inst0_O;
wire  inst1_CO;
wire  inst2_O;
wire  inst3_CO;
wire  inst4_O;
wire  inst5_CO;
wire  inst6_O;
wire  inst7_CO;
wire  inst8_O;
wire  inst9_CO;
SB_LUT4 #(.LUT_INIT(16'hC33C)) inst0 (.I0(1'b0), .I1(I0[0]), .I2(I1[0]), .I3(CIN), .O(inst0_O));
SB_CARRY inst1 (.I0(I0[0]), .I1(I1[0]), .CI(CIN), .CO(inst1_CO));
SB_LUT4 #(.LUT_INIT(16'hC33C)) inst2 (.I0(1'b0), .I1(I0[1]), .I2(I1[1]), .I3(inst1_CO), .O(inst2_O));
SB_CARRY inst3 (.I0(I0[1]), .I1(I1[1]), .CI(inst1_CO), .CO(inst3_CO));
SB_LUT4 #(.LUT_INIT(16'hC33C)) inst4 (.I0(1'b0), .I1(I0[2]), .I2(I1[2]), .I3(inst3_CO), .O(inst4_O));
SB_CARRY inst5 (.I0(I0[2]), .I1(I1[2]), .CI(inst3_CO), .CO(inst5_CO));
SB_LUT4 #(.LUT_INIT(16'hC33C)) inst6 (.I0(1'b0), .I1(I0[3]), .I2(I1[3]), .I3(inst5_CO), .O(inst6_O));
SB_CARRY inst7 (.I0(I0[3]), .I1(I1[3]), .CI(inst5_CO), .CO(inst7_CO));
SB_LUT4 #(.LUT_INIT(16'hC33C)) inst8 (.I0(1'b0), .I1(I0[4]), .I2(I1[4]), .I3(inst7_CO), .O(inst8_O));
SB_CARRY inst9 (.I0(I0[4]), .I1(I1[4]), .CI(inst7_CO), .CO(inst9_CO));
assign O = {inst8_O,inst6_O,inst4_O,inst2_O,inst0_O};
assign COUT = inst9_CO;
endmodule

module Register5CE (input [4:0] I, output [4:0] O, input  CLK, input  CE);
wire  inst0_Q;
wire  inst1_Q;
wire  inst2_Q;
wire  inst3_Q;
wire  inst4_Q;
SB_DFFE inst0 (.C(CLK), .E(CE), .D(I[0]), .Q(inst0_Q));
SB_DFFE inst1 (.C(CLK), .E(CE), .D(I[1]), .Q(inst1_Q));
SB_DFFE inst2 (.C(CLK), .E(CE), .D(I[2]), .Q(inst2_Q));
SB_DFFE inst3 (.C(CLK), .E(CE), .D(I[3]), .Q(inst3_Q));
SB_DFFE inst4 (.C(CLK), .E(CE), .D(I[4]), .Q(inst4_Q));
assign O = {inst4_Q,inst3_Q,inst2_Q,inst1_Q,inst0_Q};
endmodule

module UpDownCounter5CE (input  U, input  D, output [4:0] O, output  COUT, input  CLK, input  CE);
wire [4:0] inst0_O;
wire  inst0_COUT;
wire [4:0] inst1_O;
Addcincout5 inst0 (.I0(inst1_O), .I1({D,D,D,D,D}), .CIN(U), .O(inst0_O), .COUT(inst0_COUT));
Register5CE inst1 (.I(inst0_O), .O(inst1_O), .CLK(CLK), .CE(CE));
assign O = inst1_O;
assign COUT = inst0_COUT;
endmodule

module Mux2x8 (input [7:0] I0, input [7:0] I1, input  S, output [7:0] O);
wire  inst0_O;
wire  inst1_O;
wire  inst2_O;
wire  inst3_O;
wire  inst4_O;
wire  inst5_O;
wire  inst6_O;
wire  inst7_O;
SB_LUT4 #(.LUT_INIT(16'hCACA)) inst0 (.I0(I0[0]), .I1(I1[0]), .I2(S), .I3(1'b0), .O(inst0_O));
SB_LUT4 #(.LUT_INIT(16'hCACA)) inst1 (.I0(I0[1]), .I1(I1[1]), .I2(S), .I3(1'b0), .O(inst1_O));
SB_LUT4 #(.LUT_INIT(16'hCACA)) inst2 (.I0(I0[2]), .I1(I1[2]), .I2(S), .I3(1'b0), .O(inst2_O));
SB_LUT4 #(.LUT_INIT(16'hCACA)) inst3 (.I0(I0[3]), .I1(I1[3]), .I2(S), .I3(1'b0), .O(inst3_O));
SB_LUT4 #(.LUT_INIT(16'hCACA)) inst4 (.I0(I0[4]), .I1(I1[4]), .I2(S), .I3(1'b0), .O(inst4_O));
SB_LUT4 #(.LUT_INIT(16'hCACA)) inst5 (.I0(I0[5]), .I1(I1[5]), .I2(S), .I3(1'b0), .O(inst5_O));
SB_LUT4 #(.LUT_INIT(16'hCACA)) inst6 (.I0(I0[6]), .I1(I1[6]), .I2(S), .I3(1'b0), .O(inst6_O));
SB_LUT4 #(.LUT_INIT(16'hCACA)) inst7 (.I0(I0[7]), .I1(I1[7]), .I2(S), .I3(1'b0), .O(inst7_O));
assign O = {inst7_O,inst6_O,inst5_O,inst4_O,inst3_O,inst2_O,inst1_O,inst0_O};
endmodule

module Invert8 (input [7:0] I, output [7:0] O);
wire  inst0_O;
wire  inst1_O;
wire  inst2_O;
wire  inst3_O;
wire  inst4_O;
wire  inst5_O;
wire  inst6_O;
wire  inst7_O;
SB_LUT4 #(.LUT_INIT(16'h5555)) inst0 (.I0(I[0]), .I1(1'b0), .I2(1'b0), .I3(1'b0), .O(inst0_O));
SB_LUT4 #(.LUT_INIT(16'h5555)) inst1 (.I0(I[1]), .I1(1'b0), .I2(1'b0), .I3(1'b0), .O(inst1_O));
SB_LUT4 #(.LUT_INIT(16'h5555)) inst2 (.I0(I[2]), .I1(1'b0), .I2(1'b0), .I3(1'b0), .O(inst2_O));
SB_LUT4 #(.LUT_INIT(16'h5555)) inst3 (.I0(I[3]), .I1(1'b0), .I2(1'b0), .I3(1'b0), .O(inst3_O));
SB_LUT4 #(.LUT_INIT(16'h5555)) inst4 (.I0(I[4]), .I1(1'b0), .I2(1'b0), .I3(1'b0), .O(inst4_O));
SB_LUT4 #(.LUT_INIT(16'h5555)) inst5 (.I0(I[5]), .I1(1'b0), .I2(1'b0), .I3(1'b0), .O(inst5_O));
SB_LUT4 #(.LUT_INIT(16'h5555)) inst6 (.I0(I[6]), .I1(1'b0), .I2(1'b0), .I3(1'b0), .O(inst6_O));
SB_LUT4 #(.LUT_INIT(16'h5555)) inst7 (.I0(I[7]), .I1(1'b0), .I2(1'b0), .I3(1'b0), .O(inst7_O));
assign O = {inst7_O,inst6_O,inst5_O,inst4_O,inst3_O,inst2_O,inst1_O,inst0_O};
endmodule

module main (output  D5, output  D4, output  D3, output  D2, output  D1, input  CLKIN);
wire [17:0] inst0_O;
wire  inst0_COUT;
wire [26:0] inst1_O;
wire  inst1_COUT;
wire [1:0] inst2_O;
wire  inst2_COUT;
wire  inst3_O;
wire [7:0] inst4_O;
wire  inst4_COUT;
wire [4:0] inst5_O;
wire  inst5_COUT;
wire [7:0] inst6_O;
wire [7:0] inst7_O;
wire [7:0] inst8_O;
wire [7:0] inst9_O;
wire [7:0] inst10_O;
wire [7:0] inst11_O;
wire [7:0] inst12_O;
wire [7:0] inst13_O;
wire [7:0] inst14_O;
wire [7:0] inst15_O;
wire [7:0] inst16_O;
wire [7:0] inst17_O;
wire [7:0] inst18_O;
wire [7:0] inst19_O;
wire [7:0] inst20_O;
wire [7:0] inst21_O;
wire [7:0] inst22_O;
wire [7:0] inst23_O;
wire [7:0] inst24_O;
wire [7:0] inst25_O;
wire [7:0] inst26_O;
wire [7:0] inst27_O;
wire [7:0] inst28_O;
wire [7:0] inst29_O;
wire [7:0] inst30_O;
wire [7:0] inst31_O;
wire [7:0] inst32_O;
wire [7:0] inst33_O;
wire [7:0] inst34_O;
wire [7:0] inst35_O;
wire [7:0] inst36_O;
wire  inst37_O;
wire [7:0] inst38_O;
wire [7:0] inst39_O;
wire  inst39_COUT;
wire [7:0] inst40_O;
wire  inst40_COUT;
wire [4:0] inst41_O;
wire  inst41_COUT;
wire [7:0] inst42_O;
wire [7:0] inst43_O;
wire [7:0] inst44_O;
wire [7:0] inst45_O;
wire [7:0] inst46_O;
wire [7:0] inst47_O;
wire [7:0] inst48_O;
wire [7:0] inst49_O;
wire [7:0] inst50_O;
wire [7:0] inst51_O;
wire [7:0] inst52_O;
wire [7:0] inst53_O;
wire [7:0] inst54_O;
wire [7:0] inst55_O;
wire [7:0] inst56_O;
wire [7:0] inst57_O;
wire [7:0] inst58_O;
wire [7:0] inst59_O;
wire [7:0] inst60_O;
wire [7:0] inst61_O;
wire [7:0] inst62_O;
wire [7:0] inst63_O;
wire [7:0] inst64_O;
wire [7:0] inst65_O;
wire [7:0] inst66_O;
wire [7:0] inst67_O;
wire [7:0] inst68_O;
wire [7:0] inst69_O;
wire [7:0] inst70_O;
wire [7:0] inst71_O;
wire [7:0] inst72_O;
wire  inst73_O;
wire [7:0] inst74_O;
wire [7:0] inst75_O;
wire  inst75_COUT;
wire [7:0] inst76_O;
wire  inst76_COUT;
wire [4:0] inst77_O;
wire  inst77_COUT;
wire [7:0] inst78_O;
wire [7:0] inst79_O;
wire [7:0] inst80_O;
wire [7:0] inst81_O;
wire [7:0] inst82_O;
wire [7:0] inst83_O;
wire [7:0] inst84_O;
wire [7:0] inst85_O;
wire [7:0] inst86_O;
wire [7:0] inst87_O;
wire [7:0] inst88_O;
wire [7:0] inst89_O;
wire [7:0] inst90_O;
wire [7:0] inst91_O;
wire [7:0] inst92_O;
wire [7:0] inst93_O;
wire [7:0] inst94_O;
wire [7:0] inst95_O;
wire [7:0] inst96_O;
wire [7:0] inst97_O;
wire [7:0] inst98_O;
wire [7:0] inst99_O;
wire [7:0] inst100_O;
wire [7:0] inst101_O;
wire [7:0] inst102_O;
wire [7:0] inst103_O;
wire [7:0] inst104_O;
wire [7:0] inst105_O;
wire [7:0] inst106_O;
wire [7:0] inst107_O;
wire [7:0] inst108_O;
wire  inst109_O;
wire [7:0] inst110_O;
wire [7:0] inst111_O;
wire  inst111_COUT;
wire [7:0] inst112_O;
wire  inst112_COUT;
wire [4:0] inst113_O;
wire  inst113_COUT;
wire [7:0] inst114_O;
wire [7:0] inst115_O;
wire [7:0] inst116_O;
wire [7:0] inst117_O;
wire [7:0] inst118_O;
wire [7:0] inst119_O;
wire [7:0] inst120_O;
wire [7:0] inst121_O;
wire [7:0] inst122_O;
wire [7:0] inst123_O;
wire [7:0] inst124_O;
wire [7:0] inst125_O;
wire [7:0] inst126_O;
wire [7:0] inst127_O;
wire [7:0] inst128_O;
wire [7:0] inst129_O;
wire [7:0] inst130_O;
wire [7:0] inst131_O;
wire [7:0] inst132_O;
wire [7:0] inst133_O;
wire [7:0] inst134_O;
wire [7:0] inst135_O;
wire [7:0] inst136_O;
wire [7:0] inst137_O;
wire [7:0] inst138_O;
wire [7:0] inst139_O;
wire [7:0] inst140_O;
wire [7:0] inst141_O;
wire [7:0] inst142_O;
wire [7:0] inst143_O;
wire [7:0] inst144_O;
wire  inst145_O;
wire [7:0] inst146_O;
wire [7:0] inst147_O;
wire  inst147_COUT;
Counter18 inst0 (.O(inst0_O), .COUT(inst0_COUT), .CLK(CLKIN));
Counter27 inst1 (.O(inst1_O), .COUT(inst1_COUT), .CLK(CLKIN));
Counter2CE inst2 (.O(inst2_O), .COUT(inst2_COUT), .CLK(CLKIN), .CE(inst1_COUT));
SB_LUT4 #(.LUT_INIT(16'h6666)) inst3 (.I0(inst2_O[0]), .I1(1'b1), .I2(1'b0), .I3(1'b0), .O(inst3_O));
Counter8 inst4 (.O(inst4_O), .COUT(inst4_COUT), .CLK(CLKIN));
UpDownCounter5CE inst5 (.U(inst2_O[0]), .D(inst3_O), .O(inst5_O), .COUT(inst5_COUT), .CLK(CLKIN), .CE(inst0_COUT));
Mux2x8 inst6 (.I0({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}), .I1({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}), .S(inst5_O[0]), .O(inst6_O));
Mux2x8 inst7 (.I0({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1}), .I1({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1}), .S(inst5_O[0]), .O(inst7_O));
Mux2x8 inst8 (.I0({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0}), .I1({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0}), .S(inst5_O[0]), .O(inst8_O));
Mux2x8 inst9 (.I0({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1}), .I1({1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0}), .S(inst5_O[0]), .O(inst9_O));
Mux2x8 inst10 (.I0({1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0}), .I1({1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1}), .S(inst5_O[0]), .O(inst10_O));
Mux2x8 inst11 (.I0({1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1}), .I1({1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0}), .S(inst5_O[0]), .O(inst11_O));
Mux2x8 inst12 (.I0({1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0}), .I1({1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0}), .S(inst5_O[0]), .O(inst12_O));
Mux2x8 inst13 (.I0({1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1}), .I1({1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1}), .S(inst5_O[0]), .O(inst13_O));
Mux2x8 inst14 (.I0({1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0}), .I1({1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1}), .S(inst5_O[0]), .O(inst14_O));
Mux2x8 inst15 (.I0({1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1}), .I1({1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0}), .S(inst5_O[0]), .O(inst15_O));
Mux2x8 inst16 (.I0({1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0}), .I1({1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0}), .S(inst5_O[0]), .O(inst16_O));
Mux2x8 inst17 (.I0({1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1}), .I1({1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1}), .S(inst5_O[0]), .O(inst17_O));
Mux2x8 inst18 (.I0({1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0}), .I1({1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0}), .S(inst5_O[0]), .O(inst18_O));
Mux2x8 inst19 (.I0({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1}), .I1({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0}), .S(inst5_O[0]), .O(inst19_O));
Mux2x8 inst20 (.I0({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0}), .I1({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1}), .S(inst5_O[0]), .O(inst20_O));
Mux2x8 inst21 (.I0({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1}), .I1({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}), .S(inst5_O[0]), .O(inst21_O));
Mux2x8 inst22 (.I0(inst6_O), .I1(inst7_O), .S(inst5_O[1]), .O(inst22_O));
Mux2x8 inst23 (.I0(inst8_O), .I1(inst9_O), .S(inst5_O[1]), .O(inst23_O));
Mux2x8 inst24 (.I0(inst10_O), .I1(inst11_O), .S(inst5_O[1]), .O(inst24_O));
Mux2x8 inst25 (.I0(inst12_O), .I1(inst13_O), .S(inst5_O[1]), .O(inst25_O));
Mux2x8 inst26 (.I0(inst14_O), .I1(inst15_O), .S(inst5_O[1]), .O(inst26_O));
Mux2x8 inst27 (.I0(inst16_O), .I1(inst17_O), .S(inst5_O[1]), .O(inst27_O));
Mux2x8 inst28 (.I0(inst18_O), .I1(inst19_O), .S(inst5_O[1]), .O(inst28_O));
Mux2x8 inst29 (.I0(inst20_O), .I1(inst21_O), .S(inst5_O[1]), .O(inst29_O));
Mux2x8 inst30 (.I0(inst22_O), .I1(inst23_O), .S(inst5_O[2]), .O(inst30_O));
Mux2x8 inst31 (.I0(inst24_O), .I1(inst25_O), .S(inst5_O[2]), .O(inst31_O));
Mux2x8 inst32 (.I0(inst26_O), .I1(inst27_O), .S(inst5_O[2]), .O(inst32_O));
Mux2x8 inst33 (.I0(inst28_O), .I1(inst29_O), .S(inst5_O[2]), .O(inst33_O));
Mux2x8 inst34 (.I0(inst30_O), .I1(inst31_O), .S(inst5_O[3]), .O(inst34_O));
Mux2x8 inst35 (.I0(inst32_O), .I1(inst33_O), .S(inst5_O[3]), .O(inst35_O));
Mux2x8 inst36 (.I0(inst34_O), .I1(inst35_O), .S(inst5_O[4]), .O(inst36_O));
SB_LUT4 #(.LUT_INIT(16'h5555)) inst37 (.I0(inst39_COUT), .I1(1'b0), .I2(1'b0), .I3(1'b0), .O(inst37_O));
Invert8 inst38 (.I(inst36_O), .O(inst38_O));
Addcout8 inst39 (.I0(inst4_O), .I1(inst38_O), .O(inst39_O), .COUT(inst39_COUT));
Counter8 inst40 (.O(inst40_O), .COUT(inst40_COUT), .CLK(CLKIN));
UpDownCounter5CE inst41 (.U(inst2_O[0]), .D(inst3_O), .O(inst41_O), .COUT(inst41_COUT), .CLK(CLKIN), .CE(inst0_COUT));
Mux2x8 inst42 (.I0({1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0}), .I1({1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1}), .S(inst41_O[0]), .O(inst42_O));
Mux2x8 inst43 (.I0({1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1}), .I1({1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0}), .S(inst41_O[0]), .O(inst43_O));
Mux2x8 inst44 (.I0({1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0}), .I1({1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0}), .S(inst41_O[0]), .O(inst44_O));
Mux2x8 inst45 (.I0({1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1}), .I1({1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1}), .S(inst41_O[0]), .O(inst45_O));
Mux2x8 inst46 (.I0({1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0}), .I1({1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0}), .S(inst41_O[0]), .O(inst46_O));
Mux2x8 inst47 (.I0({1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0}), .I1({1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0}), .S(inst41_O[0]), .O(inst47_O));
Mux2x8 inst48 (.I0({1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1}), .I1({1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1}), .S(inst41_O[0]), .O(inst48_O));
Mux2x8 inst49 (.I0({1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1}), .I1({1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1}), .S(inst41_O[0]), .O(inst49_O));
Mux2x8 inst50 (.I0({1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0}), .I1({1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0}), .S(inst41_O[0]), .O(inst50_O));
Mux2x8 inst51 (.I0({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1}), .I1({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0}), .S(inst41_O[0]), .O(inst51_O));
Mux2x8 inst52 (.I0({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0}), .I1({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1}), .S(inst41_O[0]), .O(inst52_O));
Mux2x8 inst53 (.I0({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1}), .I1({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}), .S(inst41_O[0]), .O(inst53_O));
Mux2x8 inst54 (.I0({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}), .I1({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}), .S(inst41_O[0]), .O(inst54_O));
Mux2x8 inst55 (.I0({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1}), .I1({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1}), .S(inst41_O[0]), .O(inst55_O));
Mux2x8 inst56 (.I0({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0}), .I1({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0}), .S(inst41_O[0]), .O(inst56_O));
Mux2x8 inst57 (.I0({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1}), .I1({1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0}), .S(inst41_O[0]), .O(inst57_O));
Mux2x8 inst58 (.I0(inst42_O), .I1(inst43_O), .S(inst41_O[1]), .O(inst58_O));
Mux2x8 inst59 (.I0(inst44_O), .I1(inst45_O), .S(inst41_O[1]), .O(inst59_O));
Mux2x8 inst60 (.I0(inst46_O), .I1(inst47_O), .S(inst41_O[1]), .O(inst60_O));
Mux2x8 inst61 (.I0(inst48_O), .I1(inst49_O), .S(inst41_O[1]), .O(inst61_O));
Mux2x8 inst62 (.I0(inst50_O), .I1(inst51_O), .S(inst41_O[1]), .O(inst62_O));
Mux2x8 inst63 (.I0(inst52_O), .I1(inst53_O), .S(inst41_O[1]), .O(inst63_O));
Mux2x8 inst64 (.I0(inst54_O), .I1(inst55_O), .S(inst41_O[1]), .O(inst64_O));
Mux2x8 inst65 (.I0(inst56_O), .I1(inst57_O), .S(inst41_O[1]), .O(inst65_O));
Mux2x8 inst66 (.I0(inst58_O), .I1(inst59_O), .S(inst41_O[2]), .O(inst66_O));
Mux2x8 inst67 (.I0(inst60_O), .I1(inst61_O), .S(inst41_O[2]), .O(inst67_O));
Mux2x8 inst68 (.I0(inst62_O), .I1(inst63_O), .S(inst41_O[2]), .O(inst68_O));
Mux2x8 inst69 (.I0(inst64_O), .I1(inst65_O), .S(inst41_O[2]), .O(inst69_O));
Mux2x8 inst70 (.I0(inst66_O), .I1(inst67_O), .S(inst41_O[3]), .O(inst70_O));
Mux2x8 inst71 (.I0(inst68_O), .I1(inst69_O), .S(inst41_O[3]), .O(inst71_O));
Mux2x8 inst72 (.I0(inst70_O), .I1(inst71_O), .S(inst41_O[4]), .O(inst72_O));
SB_LUT4 #(.LUT_INIT(16'h5555)) inst73 (.I0(inst75_COUT), .I1(1'b0), .I2(1'b0), .I3(1'b0), .O(inst73_O));
Invert8 inst74 (.I(inst72_O), .O(inst74_O));
Addcout8 inst75 (.I0(inst40_O), .I1(inst74_O), .O(inst75_O), .COUT(inst75_COUT));
Counter8 inst76 (.O(inst76_O), .COUT(inst76_COUT), .CLK(CLKIN));
UpDownCounter5CE inst77 (.U(inst2_O[0]), .D(inst3_O), .O(inst77_O), .COUT(inst77_COUT), .CLK(CLKIN), .CE(inst0_COUT));
Mux2x8 inst78 (.I0({1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0}), .I1({1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0}), .S(inst77_O[0]), .O(inst78_O));
Mux2x8 inst79 (.I0({1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0}), .I1({1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0}), .S(inst77_O[0]), .O(inst79_O));
Mux2x8 inst80 (.I0({1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1}), .I1({1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1}), .S(inst77_O[0]), .O(inst80_O));
Mux2x8 inst81 (.I0({1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1}), .I1({1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1}), .S(inst77_O[0]), .O(inst81_O));
Mux2x8 inst82 (.I0({1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1}), .I1({1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1}), .S(inst77_O[0]), .O(inst82_O));
Mux2x8 inst83 (.I0({1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1}), .I1({1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1}), .S(inst77_O[0]), .O(inst83_O));
Mux2x8 inst84 (.I0({1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1}), .I1({1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1}), .S(inst77_O[0]), .O(inst84_O));
Mux2x8 inst85 (.I0({1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1}), .I1({1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0}), .S(inst77_O[0]), .O(inst85_O));
Mux2x8 inst86 (.I0({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}), .I1({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}), .S(inst77_O[0]), .O(inst86_O));
Mux2x8 inst87 (.I0({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1}), .I1({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1}), .S(inst77_O[0]), .O(inst87_O));
Mux2x8 inst88 (.I0({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0}), .I1({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0}), .S(inst77_O[0]), .O(inst88_O));
Mux2x8 inst89 (.I0({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1}), .I1({1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0}), .S(inst77_O[0]), .O(inst89_O));
Mux2x8 inst90 (.I0({1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0}), .I1({1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1}), .S(inst77_O[0]), .O(inst90_O));
Mux2x8 inst91 (.I0({1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1}), .I1({1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0}), .S(inst77_O[0]), .O(inst91_O));
Mux2x8 inst92 (.I0({1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0}), .I1({1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0}), .S(inst77_O[0]), .O(inst92_O));
Mux2x8 inst93 (.I0({1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1}), .I1({1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1}), .S(inst77_O[0]), .O(inst93_O));
Mux2x8 inst94 (.I0(inst78_O), .I1(inst79_O), .S(inst77_O[1]), .O(inst94_O));
Mux2x8 inst95 (.I0(inst80_O), .I1(inst81_O), .S(inst77_O[1]), .O(inst95_O));
Mux2x8 inst96 (.I0(inst82_O), .I1(inst83_O), .S(inst77_O[1]), .O(inst96_O));
Mux2x8 inst97 (.I0(inst84_O), .I1(inst85_O), .S(inst77_O[1]), .O(inst97_O));
Mux2x8 inst98 (.I0(inst86_O), .I1(inst87_O), .S(inst77_O[1]), .O(inst98_O));
Mux2x8 inst99 (.I0(inst88_O), .I1(inst89_O), .S(inst77_O[1]), .O(inst99_O));
Mux2x8 inst100 (.I0(inst90_O), .I1(inst91_O), .S(inst77_O[1]), .O(inst100_O));
Mux2x8 inst101 (.I0(inst92_O), .I1(inst93_O), .S(inst77_O[1]), .O(inst101_O));
Mux2x8 inst102 (.I0(inst94_O), .I1(inst95_O), .S(inst77_O[2]), .O(inst102_O));
Mux2x8 inst103 (.I0(inst96_O), .I1(inst97_O), .S(inst77_O[2]), .O(inst103_O));
Mux2x8 inst104 (.I0(inst98_O), .I1(inst99_O), .S(inst77_O[2]), .O(inst104_O));
Mux2x8 inst105 (.I0(inst100_O), .I1(inst101_O), .S(inst77_O[2]), .O(inst105_O));
Mux2x8 inst106 (.I0(inst102_O), .I1(inst103_O), .S(inst77_O[3]), .O(inst106_O));
Mux2x8 inst107 (.I0(inst104_O), .I1(inst105_O), .S(inst77_O[3]), .O(inst107_O));
Mux2x8 inst108 (.I0(inst106_O), .I1(inst107_O), .S(inst77_O[4]), .O(inst108_O));
SB_LUT4 #(.LUT_INIT(16'h5555)) inst109 (.I0(inst111_COUT), .I1(1'b0), .I2(1'b0), .I3(1'b0), .O(inst109_O));
Invert8 inst110 (.I(inst108_O), .O(inst110_O));
Addcout8 inst111 (.I0(inst76_O), .I1(inst110_O), .O(inst111_O), .COUT(inst111_COUT));
Counter8 inst112 (.O(inst112_O), .COUT(inst112_COUT), .CLK(CLKIN));
UpDownCounter5CE inst113 (.U(inst2_O[0]), .D(inst3_O), .O(inst113_O), .COUT(inst113_COUT), .CLK(CLKIN), .CE(inst0_COUT));
Mux2x8 inst114 (.I0({1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0}), .I1({1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1}), .S(inst113_O[0]), .O(inst114_O));
Mux2x8 inst115 (.I0({1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1}), .I1({1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1}), .S(inst113_O[0]), .O(inst115_O));
Mux2x8 inst116 (.I0({1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1}), .I1({1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1}), .S(inst113_O[0]), .O(inst116_O));
Mux2x8 inst117 (.I0({1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1}), .I1({1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1}), .S(inst113_O[0]), .O(inst117_O));
Mux2x8 inst118 (.I0({1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1}), .I1({1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1}), .S(inst113_O[0]), .O(inst118_O));
Mux2x8 inst119 (.I0({1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1}), .I1({1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b1}), .S(inst113_O[0]), .O(inst119_O));
Mux2x8 inst120 (.I0({1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0}), .I1({1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0}), .S(inst113_O[0]), .O(inst120_O));
Mux2x8 inst121 (.I0({1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0}), .I1({1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0}), .S(inst113_O[0]), .O(inst121_O));
Mux2x8 inst122 (.I0({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1}), .I1({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0}), .S(inst113_O[0]), .O(inst122_O));
Mux2x8 inst123 (.I0({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0}), .I1({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1}), .S(inst113_O[0]), .O(inst123_O));
Mux2x8 inst124 (.I0({1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0}), .I1({1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0}), .S(inst113_O[0]), .O(inst124_O));
Mux2x8 inst125 (.I0({1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1}), .I1({1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b1}), .S(inst113_O[0]), .O(inst125_O));
Mux2x8 inst126 (.I0({1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0}), .I1({1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0}), .S(inst113_O[0]), .O(inst126_O));
Mux2x8 inst127 (.I0({1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b0}), .I1({1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1}), .S(inst113_O[0]), .O(inst127_O));
Mux2x8 inst128 (.I0({1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1}), .I1({1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0}), .S(inst113_O[0]), .O(inst128_O));
Mux2x8 inst129 (.I0({1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0}), .I1({1'b0,1'b0,1'b0,1'b0,1'b1,1'b0,1'b0,1'b0}), .S(inst113_O[0]), .O(inst129_O));
Mux2x8 inst130 (.I0(inst114_O), .I1(inst115_O), .S(inst113_O[1]), .O(inst130_O));
Mux2x8 inst131 (.I0(inst116_O), .I1(inst117_O), .S(inst113_O[1]), .O(inst131_O));
Mux2x8 inst132 (.I0(inst118_O), .I1(inst119_O), .S(inst113_O[1]), .O(inst132_O));
Mux2x8 inst133 (.I0(inst120_O), .I1(inst121_O), .S(inst113_O[1]), .O(inst133_O));
Mux2x8 inst134 (.I0(inst122_O), .I1(inst123_O), .S(inst113_O[1]), .O(inst134_O));
Mux2x8 inst135 (.I0(inst124_O), .I1(inst125_O), .S(inst113_O[1]), .O(inst135_O));
Mux2x8 inst136 (.I0(inst126_O), .I1(inst127_O), .S(inst113_O[1]), .O(inst136_O));
Mux2x8 inst137 (.I0(inst128_O), .I1(inst129_O), .S(inst113_O[1]), .O(inst137_O));
Mux2x8 inst138 (.I0(inst130_O), .I1(inst131_O), .S(inst113_O[2]), .O(inst138_O));
Mux2x8 inst139 (.I0(inst132_O), .I1(inst133_O), .S(inst113_O[2]), .O(inst139_O));
Mux2x8 inst140 (.I0(inst134_O), .I1(inst135_O), .S(inst113_O[2]), .O(inst140_O));
Mux2x8 inst141 (.I0(inst136_O), .I1(inst137_O), .S(inst113_O[2]), .O(inst141_O));
Mux2x8 inst142 (.I0(inst138_O), .I1(inst139_O), .S(inst113_O[3]), .O(inst142_O));
Mux2x8 inst143 (.I0(inst140_O), .I1(inst141_O), .S(inst113_O[3]), .O(inst143_O));
Mux2x8 inst144 (.I0(inst142_O), .I1(inst143_O), .S(inst113_O[4]), .O(inst144_O));
SB_LUT4 #(.LUT_INIT(16'h5555)) inst145 (.I0(inst147_COUT), .I1(1'b0), .I2(1'b0), .I3(1'b0), .O(inst145_O));
Invert8 inst146 (.I(inst144_O), .O(inst146_O));
Addcout8 inst147 (.I0(inst112_O), .I1(inst146_O), .O(inst147_O), .COUT(inst147_COUT));
assign D5 = inst2_O[0];
assign D4 = inst145_O;
assign D3 = inst109_O;
assign D2 = inst73_O;
assign D1 = inst37_O;
endmodule

